module lab2a_circuita( 
input [2:0] v,
output [2:0] aout
);
	
assign aout = v - 3'b010;

endmodule
