module lab2a_d0(
    input [3:0] m,
    output reg [7:0] d0
);

always @(*) begin
    case(m)
        4'b0000 : d0 = 8'b11000000;
        4'b0001 : d0 = 8'b11111001;
        4'b0010 : d0 = 8'b10100100;
        4'b0011 : d0 = 8'b10110000;
        4'b0100 : d0 = 8'b10011001;
        4'b0101 : d0 = 8'b10010010;
        4'b0110 : d0 = 8'b10000010;
        4'b0111 : d0 = 8'b11111000;
        4'b1000 : d0 = 8'b10000000;
        4'b1001 : d0 = 8'b10011000;
        default : d0 = 8'b11111111;
    endcase
end

endmodule
